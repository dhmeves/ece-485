library IEEE;
use ieee.std_logic_1164.all;

entity test_bench_multicycle_datapath is
end test_bench_multicycle_datapath;

architecture behav of test_bench_multicycle_datapath is