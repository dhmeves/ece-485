library IEEE;
use ieee.std_logic_1164.all;

entity B is
	port(
		B32 : in std_logic_vector(31 downto 0);
		clk, rst, pre, ce, binvert : in std_logic;
		output : out std_logic_vector(31 downto 0)
	);
end B;

architecture behav of B is
	signal bout, b2comp : std_logic_vector(31 downto 0);
	begin
		process(clk) is
		begin 
			if rising_edge(clk) then
			if (B32(0)='1') then
				b2comp(0) <= B32(0);
				b2comp(1) <= not B32(1);
				b2comp(2) <= not B32(2);
				b2comp(3) <= not B32(3);
				b2comp(4) <= not B32(4);
				b2comp(5) <= not B32(5);
				b2comp(6) <= not B32(6);
				b2comp(7) <= not B32(7);
				b2comp(8) <= not B32(8);
				b2comp(9) <= not B32(9);
				b2comp(10) <= not B32(10);
				b2comp(11) <= not B32(11);
				b2comp(12) <= not B32(12);
				b2comp(13) <= not B32(13);
				b2comp(14) <= not B32(14);
				b2comp(15) <= not B32(15);
				b2comp(16) <= not B32(16);
				b2comp(17) <= not B32(17);
				b2comp(18) <= not B32(18);
				b2comp(19) <= not B32(19);
				b2comp(20) <= not B32(20);
				b2comp(21) <= not B32(21);
				b2comp(22) <= not B32(22);
				b2comp(23) <= not B32(23);
				b2comp(24) <= not B32(24);
				b2comp(25) <= not B32(25);
				b2comp(26) <= not B32(26);
				b2comp(27) <= not B32(27);
				b2comp(28) <= not B32(28);
				b2comp(29) <= not B32(29);
				b2comp(30) <= not B32(30);
				b2comp(31) <= not B32(31);
			elsif (B32(1)='1') then
				b2comp(0) <= B32(0);
				b2comp(1) <= B32(1);
				b2comp(2) <= not B32(2);
				b2comp(3) <= not B32(3);
				b2comp(4) <= not B32(4);
				b2comp(5) <= not B32(5);
				b2comp(6) <= not B32(6);
				b2comp(7) <= not B32(7);
				b2comp(8) <= not B32(8);
				b2comp(9) <= not B32(9);
				b2comp(10) <= not B32(10);
				b2comp(11) <= not B32(11);
				b2comp(12) <= not B32(12);
				b2comp(13) <= not B32(13);
				b2comp(14) <= not B32(14);
				b2comp(15) <= not B32(15);
				b2comp(16) <= not B32(16);
				b2comp(17) <= not B32(17);
				b2comp(18) <= not B32(18);
				b2comp(19) <= not B32(19);
				b2comp(20) <= not B32(20);
				b2comp(21) <= not B32(21);
				b2comp(22) <= not B32(22);
				b2comp(23) <= not B32(23);
				b2comp(24) <= not B32(24);
				b2comp(25) <= not B32(25);
				b2comp(26) <= not B32(26);
				b2comp(27) <= not B32(27);
				b2comp(28) <= not B32(28);
				b2comp(29) <= not B32(29);
				b2comp(30) <= not B32(30);
				b2comp(31) <= not B32(31);
			elsif (B32(2)='1') then
				b2comp(0) <= B32(0);
				b2comp(1) <= B32(1);
				b2comp(2) <= B32(2);
				b2comp(3) <= not B32(3);
				b2comp(4) <= not B32(4);
				b2comp(5) <= not B32(5);
				b2comp(6) <= not B32(6);
				b2comp(7) <= not B32(7);
				b2comp(8) <= not B32(8);
				b2comp(9) <= not B32(9);
				b2comp(10) <= not B32(10);
				b2comp(11) <= not B32(11);
				b2comp(12) <= not B32(12);
				b2comp(13) <= not B32(13);
				b2comp(14) <= not B32(14);
				b2comp(15) <= not B32(15);
				b2comp(16) <= not B32(16);
				b2comp(17) <= not B32(17);
				b2comp(18) <= not B32(18);
				b2comp(19) <= not B32(19);
				b2comp(20) <= not B32(20);
				b2comp(21) <= not B32(21);
				b2comp(22) <= not B32(22);
				b2comp(23) <= not B32(23);
				b2comp(24) <= not B32(24);
				b2comp(25) <= not B32(25);
				b2comp(26) <= not B32(26);
				b2comp(27) <= not B32(27);
				b2comp(28) <= not B32(28);
				b2comp(29) <= not B32(29);
				b2comp(30) <= not B32(30);
				b2comp(31) <= not B32(31);
			elsif (B32(3)='1') then
				b2comp(0) <= B32(0);
				b2comp(1) <= B32(1);
				b2comp(2) <= B32(2);
				b2comp(3) <= B32(3);
				b2comp(4) <= not B32(4);
				b2comp(5) <= not B32(5);
				b2comp(6) <= not B32(6);
				b2comp(7) <= not B32(7);
				b2comp(8) <= not B32(8);
				b2comp(9) <= not B32(9);
				b2comp(10) <= not B32(10);
				b2comp(11) <= not B32(11);
				b2comp(12) <= not B32(12);
				b2comp(13) <= not B32(13);
				b2comp(14) <= not B32(14);
				b2comp(15) <= not B32(15);
				b2comp(16) <= not B32(16);
				b2comp(17) <= not B32(17);
				b2comp(18) <= not B32(18);
				b2comp(19) <= not B32(19);
				b2comp(20) <= not B32(20);
				b2comp(21) <= not B32(21);
				b2comp(22) <= not B32(22);
				b2comp(23) <= not B32(23);
				b2comp(24) <= not B32(24);
				b2comp(25) <= not B32(25);
				b2comp(26) <= not B32(26);
				b2comp(27) <= not B32(27);
				b2comp(28) <= not B32(28);
				b2comp(29) <= not B32(29);
				b2comp(30) <= not B32(30);
				b2comp(31) <= not B32(31);
			elsif (B32(4)='1') then
				b2comp(0) <= B32(0);
				b2comp(1) <= B32(1);
				b2comp(2) <= B32(2);
				b2comp(3) <= B32(3);
				b2comp(4) <= B32(4);
				b2comp(5) <= not B32(5);
				b2comp(6) <= not B32(6);
				b2comp(7) <= not B32(7);
				b2comp(8) <= not B32(8);
				b2comp(9) <= not B32(9);
				b2comp(10) <= not B32(10);
				b2comp(11) <= not B32(11);
				b2comp(12) <= not B32(12);
				b2comp(13) <= not B32(13);
				b2comp(14) <= not B32(14);
				b2comp(15) <= not B32(15);
				b2comp(16) <= not B32(16);
				b2comp(17) <= not B32(17);
				b2comp(18) <= not B32(18);
				b2comp(19) <= not B32(19);
				b2comp(20) <= not B32(20);
				b2comp(21) <= not B32(21);
				b2comp(22) <= not B32(22);
				b2comp(23) <= not B32(23);
				b2comp(24) <= not B32(24);
				b2comp(25) <= not B32(25);
				b2comp(26) <= not B32(26);
				b2comp(27) <= not B32(27);
				b2comp(28) <= not B32(28);
				b2comp(29) <= not B32(29);
				b2comp(30) <= not B32(30);
				b2comp(31) <= not B32(31);
			elsif (B32(5)='1') then
				b2comp(0) <= B32(0);
				b2comp(1) <= B32(1);
				b2comp(2) <= B32(2);
				b2comp(3) <= B32(3);
				b2comp(4) <= B32(4);
				b2comp(5) <= B32(5);
				b2comp(6) <= not B32(6);
				b2comp(7) <= not B32(7);
				b2comp(8) <= not B32(8);
				b2comp(9) <= not B32(9);
				b2comp(10) <= not B32(10);
				b2comp(11) <= not B32(11);
				b2comp(12) <= not B32(12);
				b2comp(13) <= not B32(13);
				b2comp(14) <= not B32(14);
				b2comp(15) <= not B32(15);
				b2comp(16) <= not B32(16);
				b2comp(17) <= not B32(17);
				b2comp(18) <= not B32(18);
				b2comp(19) <= not B32(19);
				b2comp(20) <= not B32(20);
				b2comp(21) <= not B32(21);
				b2comp(22) <= not B32(22);
				b2comp(23) <= not B32(23);
				b2comp(24) <= not B32(24);
				b2comp(25) <= not B32(25);
				b2comp(26) <= not B32(26);
				b2comp(27) <= not B32(27);
				b2comp(28) <= not B32(28);
				b2comp(29) <= not B32(29);
				b2comp(30) <= not B32(30);
				b2comp(31) <= not B32(31);
			elsif (B32(6)='1') then
				b2comp(0) <= B32(0);
				b2comp(1) <= B32(1);
				b2comp(2) <= B32(2);
				b2comp(3) <= B32(3);
				b2comp(4) <= B32(4);
				b2comp(5) <= B32(5);
				b2comp(6) <= B32(6);
				b2comp(7) <= not B32(7);
				b2comp(8) <= not B32(8);
				b2comp(9) <= not B32(9);
				b2comp(10) <= not B32(10);
				b2comp(11) <= not B32(11);
				b2comp(12) <= not B32(12);
				b2comp(13) <= not B32(13);
				b2comp(14) <= not B32(14);
				b2comp(15) <= not B32(15);
				b2comp(16) <= not B32(16);
				b2comp(17) <= not B32(17);
				b2comp(18) <= not B32(18);
				b2comp(19) <= not B32(19);
				b2comp(20) <= not B32(20);
				b2comp(21) <= not B32(21);
				b2comp(22) <= not B32(22);
				b2comp(23) <= not B32(23);
				b2comp(24) <= not B32(24);
				b2comp(25) <= not B32(25);
				b2comp(26) <= not B32(26);
				b2comp(27) <= not B32(27);
				b2comp(28) <= not B32(28);
				b2comp(29) <= not B32(29);
				b2comp(30) <= not B32(30);
				b2comp(31) <= not B32(31);
			elsif (B32(7)='1') then
				b2comp(0) <= B32(0);
				b2comp(1) <= B32(1);
				b2comp(2) <= B32(2);
				b2comp(3) <= B32(3);
				b2comp(4) <= B32(4);
				b2comp(5) <= B32(5);
				b2comp(6) <= B32(6);
				b2comp(7) <= B32(7);
				b2comp(8) <= not B32(8);
				b2comp(9) <= not B32(9);
				b2comp(10) <= not B32(10);
				b2comp(11) <= not B32(11);
				b2comp(12) <= not B32(12);
				b2comp(13) <= not B32(13);
				b2comp(14) <= not B32(14);
				b2comp(15) <= not B32(15);
				b2comp(16) <= not B32(16);
				b2comp(17) <= not B32(17);
				b2comp(18) <= not B32(18);
				b2comp(19) <= not B32(19);
				b2comp(20) <= not B32(20);
				b2comp(21) <= not B32(21);
				b2comp(22) <= not B32(22);
				b2comp(23) <= not B32(23);
				b2comp(24) <= not B32(24);
				b2comp(25) <= not B32(25);
				b2comp(26) <= not B32(26);
				b2comp(27) <= not B32(27);
				b2comp(28) <= not B32(28);
				b2comp(29) <= not B32(29);
				b2comp(30) <= not B32(30);
				b2comp(31) <= not B32(31);
			elsif (B32(8)='1') then
				b2comp(0) <= B32(0);
				b2comp(1) <= B32(1);
				b2comp(2) <= B32(2);
				b2comp(3) <= B32(3);
				b2comp(4) <= B32(4);
				b2comp(5) <= B32(5);
				b2comp(6) <= B32(6);
				b2comp(7) <= B32(7);
				b2comp(8) <= B32(8);
				b2comp(9) <= not B32(9);
				b2comp(10) <= not B32(10);
				b2comp(11) <= not B32(11);
				b2comp(12) <= not B32(12);
				b2comp(13) <= not B32(13);
				b2comp(14) <= not B32(14);
				b2comp(15) <= not B32(15);
				b2comp(16) <= not B32(16);
				b2comp(17) <= not B32(17);
				b2comp(18) <= not B32(18);
				b2comp(19) <= not B32(19);
				b2comp(20) <= not B32(20);
				b2comp(21) <= not B32(21);
				b2comp(22) <= not B32(22);
				b2comp(23) <= not B32(23);
				b2comp(24) <= not B32(24);
				b2comp(25) <= not B32(25);
				b2comp(26) <= not B32(26);
				b2comp(27) <= not B32(27);
				b2comp(28) <= not B32(28);
				b2comp(29) <= not B32(29);
				b2comp(30) <= not B32(30);
				b2comp(31) <= not B32(31);
			elsif (B32(9)='1') then
				b2comp(0) <= B32(0);
				b2comp(1) <= B32(1);
				b2comp(2) <= B32(2);
				b2comp(3) <= B32(3);
				b2comp(4) <= B32(4);
				b2comp(5) <= B32(5);
				b2comp(6) <= B32(6);
				b2comp(7) <= B32(7);
				b2comp(8) <= B32(8);
				b2comp(9) <= B32(9);
				b2comp(10) <= not B32(10);
				b2comp(11) <= not B32(11);
				b2comp(12) <= not B32(12);
				b2comp(13) <= not B32(13);
				b2comp(14) <= not B32(14);
				b2comp(15) <= not B32(15);
				b2comp(16) <= not B32(16);
				b2comp(17) <= not B32(17);
				b2comp(18) <= not B32(18);
				b2comp(19) <= not B32(19);
				b2comp(20) <= not B32(20);
				b2comp(21) <= not B32(21);
				b2comp(22) <= not B32(22);
				b2comp(23) <= not B32(23);
				b2comp(24) <= not B32(24);
				b2comp(25) <= not B32(25);
				b2comp(26) <= not B32(26);
				b2comp(27) <= not B32(27);
				b2comp(28) <= not B32(28);
				b2comp(29) <= not B32(29);
				b2comp(30) <= not B32(30);
				b2comp(31) <= not B32(31);
			elsif (B32(10)='1') then
				b2comp(0) <= B32(0);
				b2comp(1) <= B32(1);
				b2comp(2) <= B32(2);
				b2comp(3) <= B32(3);
				b2comp(4) <= B32(4);
				b2comp(5) <= B32(5);
				b2comp(6) <= B32(6);
				b2comp(7) <= B32(7);
				b2comp(8) <= B32(8);
				b2comp(9) <= B32(9);
				b2comp(10) <= B32(10);
				b2comp(11) <= not B32(11);
				b2comp(12) <= not B32(12);
				b2comp(13) <= not B32(13);
				b2comp(14) <= not B32(14);
				b2comp(15) <= not B32(15);
				b2comp(16) <= not B32(16);
				b2comp(17) <= not B32(17);
				b2comp(18) <= not B32(18);
				b2comp(19) <= not B32(19);
				b2comp(20) <= not B32(20);
				b2comp(21) <= not B32(21);
				b2comp(22) <= not B32(22);
				b2comp(23) <= not B32(23);
				b2comp(24) <= not B32(24);
				b2comp(25) <= not B32(25);
				b2comp(26) <= not B32(26);
				b2comp(27) <= not B32(27);
				b2comp(28) <= not B32(28);
				b2comp(29) <= not B32(29);
				b2comp(30) <= not B32(30);
				b2comp(31) <= not B32(31);
			elsif (B32(11)='1') then
				b2comp(0) <= B32(0);
				b2comp(1) <= B32(1);
				b2comp(2) <= B32(2);
				b2comp(3) <= B32(3);
				b2comp(4) <= B32(4);
				b2comp(5) <= B32(5);
				b2comp(6) <= B32(6);
				b2comp(7) <= B32(7);
				b2comp(8) <= B32(8);
				b2comp(9) <= B32(9);
				b2comp(10) <= B32(10);
				b2comp(11) <= B32(11);
				b2comp(12) <= not B32(12);
				b2comp(13) <= not B32(13);
				b2comp(14) <= not B32(14);
				b2comp(15) <= not B32(15);
				b2comp(16) <= not B32(16);
				b2comp(17) <= not B32(17);
				b2comp(18) <= not B32(18);
				b2comp(19) <= not B32(19);
				b2comp(20) <= not B32(20);
				b2comp(21) <= not B32(21);
				b2comp(22) <= not B32(22);
				b2comp(23) <= not B32(23);
				b2comp(24) <= not B32(24);
				b2comp(25) <= not B32(25);
				b2comp(26) <= not B32(26);
				b2comp(27) <= not B32(27);
				b2comp(28) <= not B32(28);
				b2comp(29) <= not B32(29);
				b2comp(30) <= not B32(30);
				b2comp(31) <= not B32(31);
			elsif (B32(12)='1') then
				b2comp(0) <= B32(0);
				b2comp(1) <= B32(1);
				b2comp(2) <= B32(2);
				b2comp(3) <= B32(3);
				b2comp(4) <= B32(4);
				b2comp(5) <= B32(5);
				b2comp(6) <= B32(6);
				b2comp(7) <= B32(7);
				b2comp(8) <= B32(8);
				b2comp(9) <= B32(9);
				b2comp(10) <= B32(10);
				b2comp(11) <= B32(11);
				b2comp(12) <= B32(12);
				b2comp(13) <= not B32(13);
				b2comp(14) <= not B32(14);
				b2comp(15) <= not B32(15);
				b2comp(16) <= not B32(16);
				b2comp(17) <= not B32(17);
				b2comp(18) <= not B32(18);
				b2comp(19) <= not B32(19);
				b2comp(20) <= not B32(20);
				b2comp(21) <= not B32(21);
				b2comp(22) <= not B32(22);
				b2comp(23) <= not B32(23);
				b2comp(24) <= not B32(24);
				b2comp(25) <= not B32(25);
				b2comp(26) <= not B32(26);
				b2comp(27) <= not B32(27);
				b2comp(28) <= not B32(28);
				b2comp(29) <= not B32(29);
				b2comp(30) <= not B32(30);
				b2comp(31) <= not B32(31);
			elsif (B32(13)='1') then
				b2comp(0) <= B32(0);
				b2comp(1) <= B32(1);
				b2comp(2) <= B32(2);
				b2comp(3) <= B32(3);
				b2comp(4) <= B32(4);
				b2comp(5) <= B32(5);
				b2comp(6) <= B32(6);
				b2comp(7) <= B32(7);
				b2comp(8) <= B32(8);
				b2comp(9) <= B32(9);
				b2comp(10) <= B32(10);
				b2comp(11) <= B32(11);
				b2comp(12) <= B32(12);
				b2comp(13) <= B32(13);
				b2comp(14) <= not B32(14);
				b2comp(15) <= not B32(15);
				b2comp(16) <= not B32(16);
				b2comp(17) <= not B32(17);
				b2comp(18) <= not B32(18);
				b2comp(19) <= not B32(19);
				b2comp(20) <= not B32(20);
				b2comp(21) <= not B32(21);
				b2comp(22) <= not B32(22);
				b2comp(23) <= not B32(23);
				b2comp(24) <= not B32(24);
				b2comp(25) <= not B32(25);
				b2comp(26) <= not B32(26);
				b2comp(27) <= not B32(27);
				b2comp(28) <= not B32(28);
				b2comp(29) <= not B32(29);
				b2comp(30) <= not B32(30);
				b2comp(31) <= not B32(31);
			elsif (B32(14)='1') then
				b2comp(0) <= B32(0);
				b2comp(1) <= B32(1);
				b2comp(2) <= B32(2);
				b2comp(3) <= B32(3);
				b2comp(4) <= B32(4);
				b2comp(5) <= B32(5);
				b2comp(6) <= B32(6);
				b2comp(7) <= B32(7);
				b2comp(8) <= B32(8);
				b2comp(9) <= B32(9);
				b2comp(10) <= B32(10);
				b2comp(11) <= B32(11);
				b2comp(12) <= B32(12);
				b2comp(13) <= B32(13);
				b2comp(14) <= B32(14);
				b2comp(15) <= not B32(15);
				b2comp(16) <= not B32(16);
				b2comp(17) <= not B32(17);
				b2comp(18) <= not B32(18);
				b2comp(19) <= not B32(19);
				b2comp(20) <= not B32(20);
				b2comp(21) <= not B32(21);
				b2comp(22) <= not B32(22);
				b2comp(23) <= not B32(23);
				b2comp(24) <= not B32(24);
				b2comp(25) <= not B32(25);
				b2comp(26) <= not B32(26);
				b2comp(27) <= not B32(27);
				b2comp(28) <= not B32(28);
				b2comp(29) <= not B32(29);
				b2comp(30) <= not B32(30);
				b2comp(31) <= not B32(31);
			elsif (B32(15)='1') then
				b2comp(0) <= B32(0);
				b2comp(1) <= B32(1);
				b2comp(2) <= B32(2);
				b2comp(3) <= B32(3);
				b2comp(4) <= B32(4);
				b2comp(5) <= B32(5);
				b2comp(6) <= B32(6);
				b2comp(7) <= B32(7);
				b2comp(8) <= B32(8);
				b2comp(9) <= B32(9);
				b2comp(10) <= B32(10);
				b2comp(11) <= B32(11);
				b2comp(12) <= B32(12);
				b2comp(13) <= B32(13);
				b2comp(14) <= B32(14);
				b2comp(15) <= B32(15);
				b2comp(16) <= not B32(16);
				b2comp(17) <= not B32(17);
				b2comp(18) <= not B32(18);
				b2comp(19) <= not B32(19);
				b2comp(20) <= not B32(20);
				b2comp(21) <= not B32(21);
				b2comp(22) <= not B32(22);
				b2comp(23) <= not B32(23);
				b2comp(24) <= not B32(24);
				b2comp(25) <= not B32(25);
				b2comp(26) <= not B32(26);
				b2comp(27) <= not B32(27);
				b2comp(28) <= not B32(28);
				b2comp(29) <= not B32(29);
				b2comp(30) <= not B32(30);
				b2comp(31) <= not B32(31);
			elsif (B32(16)='1') then
				b2comp(0) <= B32(0);
				b2comp(1) <= B32(1);
				b2comp(2) <= B32(2);
				b2comp(3) <= B32(3);
				b2comp(4) <= B32(4);
				b2comp(5) <= B32(5);
				b2comp(6) <= B32(6);
				b2comp(7) <= B32(7);
				b2comp(8) <= B32(8);
				b2comp(9) <= B32(9);
				b2comp(10) <= B32(10);
				b2comp(11) <= B32(11);
				b2comp(12) <= B32(12);
				b2comp(13) <= B32(13);
				b2comp(14) <= B32(14);
				b2comp(15) <= B32(15);
				b2comp(16) <= B32(16);
				b2comp(17) <= not B32(17);
				b2comp(18) <= not B32(18);
				b2comp(19) <= not B32(19);
				b2comp(20) <= not B32(20);
				b2comp(21) <= not B32(21);
				b2comp(22) <= not B32(22);
				b2comp(23) <= not B32(23);
				b2comp(24) <= not B32(24);
				b2comp(25) <= not B32(25);
				b2comp(26) <= not B32(26);
				b2comp(27) <= not B32(27);
				b2comp(28) <= not B32(28);
				b2comp(29) <= not B32(29);
				b2comp(30) <= not B32(30);
				b2comp(31) <= not B32(31);
			elsif (B32(17)='1') then
				b2comp(0) <= B32(0);
				b2comp(1) <= B32(1);
				b2comp(2) <= B32(2);
				b2comp(3) <= B32(3);
				b2comp(4) <= B32(4);
				b2comp(5) <= B32(5);
				b2comp(6) <= B32(6);
				b2comp(7) <= B32(7);
				b2comp(8) <= B32(8);
				b2comp(9) <= B32(9);
				b2comp(10) <= B32(10);
				b2comp(11) <= B32(11);
				b2comp(12) <= B32(12);
				b2comp(13) <= B32(13);
				b2comp(14) <= B32(14);
				b2comp(15) <= B32(15);
				b2comp(16) <= B32(16);
				b2comp(17) <= B32(17);
				b2comp(18) <= not B32(18);
				b2comp(19) <= not B32(19);
				b2comp(20) <= not B32(20);
				b2comp(21) <= not B32(21);
				b2comp(22) <= not B32(22);
				b2comp(23) <= not B32(23);
				b2comp(24) <= not B32(24);
				b2comp(25) <= not B32(25);
				b2comp(26) <= not B32(26);
				b2comp(27) <= not B32(27);
				b2comp(28) <= not B32(28);
				b2comp(29) <= not B32(29);
				b2comp(30) <= not B32(30);
				b2comp(31) <= not B32(31);
			elsif (B32(18)='1') then
				b2comp(0) <= B32(0);
				b2comp(1) <= B32(1);
				b2comp(2) <= B32(2);
				b2comp(3) <= B32(3);
				b2comp(4) <= B32(4);
				b2comp(5) <= B32(5);
				b2comp(6) <= B32(6);
				b2comp(7) <= B32(7);
				b2comp(8) <= B32(8);
				b2comp(9) <= B32(9);
				b2comp(10) <= B32(10);
				b2comp(11) <= B32(11);
				b2comp(12) <= B32(12);
				b2comp(13) <= B32(13);
				b2comp(14) <= B32(14);
				b2comp(15) <= B32(15);
				b2comp(16) <= B32(16);
				b2comp(17) <= B32(17);
				b2comp(18) <= B32(18);
				b2comp(19) <= not B32(19);
				b2comp(20) <= not B32(20);
				b2comp(21) <= not B32(21);
				b2comp(22) <= not B32(22);
				b2comp(23) <= not B32(23);
				b2comp(24) <= not B32(24);
				b2comp(25) <= not B32(25);
				b2comp(26) <= not B32(26);
				b2comp(27) <= not B32(27);
				b2comp(28) <= not B32(28);
				b2comp(29) <= not B32(29);
				b2comp(30) <= not B32(30);
				b2comp(31) <= not B32(31);
			elsif (B32(19)='1') then
				b2comp(0) <= B32(0);
				b2comp(1) <= B32(1);
				b2comp(2) <= B32(2);
				b2comp(3) <= B32(3);
				b2comp(4) <= B32(4);
				b2comp(5) <= B32(5);
				b2comp(6) <= B32(6);
				b2comp(7) <= B32(7);
				b2comp(8) <= B32(8);
				b2comp(9) <= B32(9);
				b2comp(10) <= B32(10);
				b2comp(11) <= B32(11);
				b2comp(12) <= B32(12);
				b2comp(13) <= B32(13);
				b2comp(14) <= B32(14);
				b2comp(15) <= B32(15);
				b2comp(16) <= B32(16);
				b2comp(17) <= B32(17);
				b2comp(18) <= B32(18);
				b2comp(19) <= B32(19);
				b2comp(20) <= not B32(20);
				b2comp(21) <= not B32(21);
				b2comp(22) <= not B32(22);
				b2comp(23) <= not B32(23);
				b2comp(24) <= not B32(24);
				b2comp(25) <= not B32(25);
				b2comp(26) <= not B32(26);
				b2comp(27) <= not B32(27);
				b2comp(28) <= not B32(28);
				b2comp(29) <= not B32(29);
				b2comp(30) <= not B32(30);
				b2comp(31) <= not B32(31);
			elsif (B32(20)='1') then
				b2comp(0) <= B32(0);
				b2comp(1) <= B32(1);
				b2comp(2) <= B32(2);
				b2comp(3) <= B32(3);
				b2comp(4) <= B32(4);
				b2comp(5) <= B32(5);
				b2comp(6) <= B32(6);
				b2comp(7) <= B32(7);
				b2comp(8) <= B32(8);
				b2comp(9) <= B32(9);
				b2comp(10) <= B32(10);
				b2comp(11) <= B32(11);
				b2comp(12) <= B32(12);
				b2comp(13) <= B32(13);
				b2comp(14) <= B32(14);
				b2comp(15) <= B32(15);
				b2comp(16) <= B32(16);
				b2comp(17) <= B32(17);
				b2comp(18) <= B32(18);
				b2comp(19) <= B32(19);
				b2comp(20) <= B32(20);
				b2comp(21) <= not B32(21);
				b2comp(22) <= not B32(22);
				b2comp(23) <= not B32(23);
				b2comp(24) <= not B32(24);
				b2comp(25) <= not B32(25);
				b2comp(26) <= not B32(26);
				b2comp(27) <= not B32(27);
				b2comp(28) <= not B32(28);
				b2comp(29) <= not B32(29);
				b2comp(30) <= not B32(30);
				b2comp(31) <= not B32(31);
			elsif (B32(21)='1') then
				b2comp(0) <= B32(0);
				b2comp(1) <= B32(1);
				b2comp(2) <= B32(2);
				b2comp(3) <= B32(3);
				b2comp(4) <= B32(4);
				b2comp(5) <= B32(5);
				b2comp(6) <= B32(6);
				b2comp(7) <= B32(7);
				b2comp(8) <= B32(8);
				b2comp(9) <= B32(9);
				b2comp(10) <= B32(10);
				b2comp(11) <= B32(11);
				b2comp(12) <= B32(12);
				b2comp(13) <= B32(13);
				b2comp(14) <= B32(14);
				b2comp(15) <= B32(15);
				b2comp(16) <= B32(16);
				b2comp(17) <= B32(17);
				b2comp(18) <= B32(18);
				b2comp(19) <= B32(19);
				b2comp(20) <= B32(20);
				b2comp(21) <= B32(21);
				b2comp(22) <= not B32(22);
				b2comp(23) <= not B32(23);
				b2comp(24) <= not B32(24);
				b2comp(25) <= not B32(25);
				b2comp(26) <= not B32(26);
				b2comp(27) <= not B32(27);
				b2comp(28) <= not B32(28);
				b2comp(29) <= not B32(29);
				b2comp(30) <= not B32(30);
				b2comp(31) <= not B32(31);
			elsif (B32(22)='1') then
				b2comp(0) <= B32(0);
				b2comp(1) <= B32(1);
				b2comp(2) <= B32(2);
				b2comp(3) <= B32(3);
				b2comp(4) <= B32(4);
				b2comp(5) <= B32(5);
				b2comp(6) <= B32(6);
				b2comp(7) <= B32(7);
				b2comp(8) <= B32(8);
				b2comp(9) <= B32(9);
				b2comp(10) <= B32(10);
				b2comp(11) <= B32(11);
				b2comp(12) <= B32(12);
				b2comp(13) <= B32(13);
				b2comp(14) <= B32(14);
				b2comp(15) <= B32(15);
				b2comp(16) <= B32(16);
				b2comp(17) <= B32(17);
				b2comp(18) <= B32(18);
				b2comp(19) <= B32(19);
				b2comp(20) <= B32(20);
				b2comp(21) <= B32(21);
				b2comp(22) <= B32(22);
				b2comp(23) <= not B32(23);
				b2comp(24) <= not B32(24);
				b2comp(25) <= not B32(25);
				b2comp(26) <= not B32(26);
				b2comp(27) <= not B32(27);
				b2comp(28) <= not B32(28);
				b2comp(29) <= not B32(29);
				b2comp(30) <= not B32(30);
				b2comp(31) <= not B32(31);
			elsif (B32(23)='1') then
				b2comp(0) <= B32(0);
				b2comp(1) <= B32(1);
				b2comp(2) <= B32(2);
				b2comp(3) <= B32(3);
				b2comp(4) <= B32(4);
				b2comp(5) <= B32(5);
				b2comp(6) <= B32(6);
				b2comp(7) <= B32(7);
				b2comp(8) <= B32(8);
				b2comp(9) <= B32(9);
				b2comp(10) <= B32(10);
				b2comp(11) <= B32(11);
				b2comp(12) <= B32(12);
				b2comp(13) <= B32(13);
				b2comp(14) <= B32(14);
				b2comp(15) <= B32(15);
				b2comp(16) <= B32(16);
				b2comp(17) <= B32(17);
				b2comp(18) <= B32(18);
				b2comp(19) <= B32(19);
				b2comp(20) <= B32(20);
				b2comp(21) <= B32(21);
				b2comp(22) <= B32(22);
				b2comp(23) <= B32(23);
				b2comp(24) <= not B32(24);
				b2comp(25) <= not B32(25);
				b2comp(26) <= not B32(26);
				b2comp(27) <= not B32(27);
				b2comp(28) <= not B32(28);
				b2comp(29) <= not B32(29);
				b2comp(30) <= not B32(30);
				b2comp(31) <= not B32(31);
			elsif (B32(24)='1') then
				b2comp(0) <= B32(0);
				b2comp(1) <= B32(1);
				b2comp(2) <= B32(2);
				b2comp(3) <= B32(3);
				b2comp(4) <= B32(4);
				b2comp(5) <= B32(5);
				b2comp(6) <= B32(6);
				b2comp(7) <= B32(7);
				b2comp(8) <= B32(8);
				b2comp(9) <= B32(9);
				b2comp(10) <= B32(10);
				b2comp(11) <= B32(11);
				b2comp(12) <= B32(12);
				b2comp(13) <= B32(13);
				b2comp(14) <= B32(14);
				b2comp(15) <= B32(15);
				b2comp(16) <= B32(16);
				b2comp(17) <= B32(17);
				b2comp(18) <= B32(18);
				b2comp(19) <= B32(19);
				b2comp(20) <= B32(20);
				b2comp(21) <= B32(21);
				b2comp(22) <= B32(22);
				b2comp(23) <= B32(23);
				b2comp(24) <= B32(24);
				b2comp(25) <= not B32(25);
				b2comp(26) <= not B32(26);
				b2comp(27) <= not B32(27);
				b2comp(28) <= not B32(28);
				b2comp(29) <= not B32(29);
				b2comp(30) <= not B32(30);
				b2comp(31) <= not B32(31);
			elsif (B32(25)='1') then
				b2comp(0) <= B32(0);
				b2comp(1) <= B32(1);
				b2comp(2) <= B32(2);
				b2comp(3) <= B32(3);
				b2comp(4) <= B32(4);
				b2comp(5) <= B32(5);
				b2comp(6) <= B32(6);
				b2comp(7) <= B32(7);
				b2comp(8) <= B32(8);
				b2comp(9) <= B32(9);
				b2comp(10) <= B32(10);
				b2comp(11) <= B32(11);
				b2comp(12) <= B32(12);
				b2comp(13) <= B32(13);
				b2comp(14) <= B32(14);
				b2comp(15) <= B32(15);
				b2comp(16) <= B32(16);
				b2comp(17) <= B32(17);
				b2comp(18) <= B32(18);
				b2comp(19) <= B32(19);
				b2comp(20) <= B32(20);
				b2comp(21) <= B32(21);
				b2comp(22) <= B32(22);
				b2comp(23) <= B32(23);
				b2comp(24) <= B32(24);
				b2comp(25) <= B32(25);
				b2comp(26) <= not B32(26);
				b2comp(27) <= not B32(27);
				b2comp(28) <= not B32(28);
				b2comp(29) <= not B32(29);
				b2comp(30) <= not B32(30);
				b2comp(31) <= not B32(31);
			elsif (B32(26)='1') then
				b2comp(0) <= B32(0);
				b2comp(1) <= B32(1);
				b2comp(2) <= B32(2);
				b2comp(3) <= B32(3);
				b2comp(4) <= B32(4);
				b2comp(5) <= B32(5);
				b2comp(6) <= B32(6);
				b2comp(7) <= B32(7);
				b2comp(8) <= B32(8);
				b2comp(9) <= B32(9);
				b2comp(10) <= B32(10);
				b2comp(11) <= B32(11);
				b2comp(12) <= B32(12);
				b2comp(13) <= B32(13);
				b2comp(14) <= B32(14);
				b2comp(15) <= B32(15);
				b2comp(16) <= B32(16);
				b2comp(17) <= B32(17);
				b2comp(18) <= B32(18);
				b2comp(19) <= B32(19);
				b2comp(20) <= B32(20);
				b2comp(21) <= B32(21);
				b2comp(22) <= B32(22);
				b2comp(23) <= B32(23);
				b2comp(24) <= B32(24);
				b2comp(25) <= B32(25);
				b2comp(26) <= B32(26);
				b2comp(27) <= not B32(27);
				b2comp(28) <= not B32(28);
				b2comp(29) <= not B32(29);
				b2comp(30) <= not B32(30);
				b2comp(31) <= not B32(31);
			elsif (B32(27)='1') then
				b2comp(0) <= B32(0);
				b2comp(1) <= B32(1);
				b2comp(2) <= B32(2);
				b2comp(3) <= B32(3);
				b2comp(4) <= B32(4);
				b2comp(5) <= B32(5);
				b2comp(6) <= B32(6);
				b2comp(7) <= B32(7);
				b2comp(8) <= B32(8);
				b2comp(9) <= B32(9);
				b2comp(10) <= B32(10);
				b2comp(11) <= B32(11);
				b2comp(12) <= B32(12);
				b2comp(13) <= B32(13);
				b2comp(14) <= B32(14);
				b2comp(15) <= B32(15);
				b2comp(16) <= B32(16);
				b2comp(17) <= B32(17);
				b2comp(18) <= B32(18);
				b2comp(19) <= B32(19);
				b2comp(20) <= B32(20);
				b2comp(21) <= B32(21);
				b2comp(22) <= B32(22);
				b2comp(23) <= B32(23);
				b2comp(24) <= B32(24);
				b2comp(25) <= B32(25);
				b2comp(26) <= B32(26);
				b2comp(27) <= B32(27);
				b2comp(28) <= not B32(28);
				b2comp(29) <= not B32(29);
				b2comp(30) <= not B32(30);
				b2comp(31) <= not B32(31);
			elsif (B32(28)='1') then
				b2comp(0) <= B32(0);
				b2comp(1) <= B32(1);
				b2comp(2) <= B32(2);
				b2comp(3) <= B32(3);
				b2comp(4) <= B32(4);
				b2comp(5) <= B32(5);
				b2comp(6) <= B32(6);
				b2comp(7) <= B32(7);
				b2comp(8) <= B32(8);
				b2comp(9) <= B32(9);
				b2comp(10) <= B32(10);
				b2comp(11) <= B32(11);
				b2comp(12) <= B32(12);
				b2comp(13) <= B32(13);
				b2comp(14) <= B32(14);
				b2comp(15) <= B32(15);
				b2comp(16) <= B32(16);
				b2comp(17) <= B32(17);
				b2comp(18) <= B32(18);
				b2comp(19) <= B32(19);
				b2comp(20) <= B32(20);
				b2comp(21) <= B32(21);
				b2comp(22) <= B32(22);
				b2comp(23) <= B32(23);
				b2comp(24) <= B32(24);
				b2comp(25) <= B32(25);
				b2comp(26) <= B32(26);
				b2comp(27) <= B32(27);
				b2comp(28) <= B32(28);
				b2comp(29) <= not B32(29);
				b2comp(30) <= not B32(30);
				b2comp(31) <= not B32(31);
			elsif (B32(29)='1') then
				b2comp(0) <= B32(0);
				b2comp(1) <= B32(1);
				b2comp(2) <= B32(2);
				b2comp(3) <= B32(3);
				b2comp(4) <= B32(4);
				b2comp(5) <= B32(5);
				b2comp(6) <= B32(6);
				b2comp(7) <= B32(7);
				b2comp(8) <= B32(8);
				b2comp(9) <= B32(9);
				b2comp(10) <= B32(10);
				b2comp(11) <= B32(11);
				b2comp(12) <= B32(12);
				b2comp(13) <= B32(13);
				b2comp(14) <= B32(14);
				b2comp(15) <= B32(15);
				b2comp(16) <= B32(16);
				b2comp(17) <= B32(17);
				b2comp(18) <= B32(18);
				b2comp(19) <= B32(19);
				b2comp(20) <= B32(20);
				b2comp(21) <= B32(21);
				b2comp(22) <= B32(22);
				b2comp(23) <= B32(23);
				b2comp(24) <= B32(24);
				b2comp(25) <= B32(25);
				b2comp(26) <= B32(26);
				b2comp(27) <= B32(27);
				b2comp(28) <= B32(28);
				b2comp(29) <= B32(29);
				b2comp(30) <= not B32(30);
				b2comp(31) <= not B32(31);
			elsif (B32(30)='1') then
				b2comp(0) <= B32(0);
				b2comp(1) <= B32(1);
				b2comp(2) <= B32(2);
				b2comp(3) <= B32(3);
				b2comp(4) <= B32(4);
				b2comp(5) <= B32(5);
				b2comp(6) <= B32(6);
				b2comp(7) <= B32(7);
				b2comp(8) <= B32(8);
				b2comp(9) <= B32(9);
				b2comp(10) <= B32(10);
				b2comp(11) <= B32(11);
				b2comp(12) <= B32(12);
				b2comp(13) <= B32(13);
				b2comp(14) <= B32(14);
				b2comp(15) <= B32(15);
				b2comp(16) <= B32(16);
				b2comp(17) <= B32(17);
				b2comp(18) <= B32(18);
				b2comp(19) <= B32(19);
				b2comp(20) <= B32(20);
				b2comp(21) <= B32(21);
				b2comp(22) <= B32(22);
				b2comp(23) <= B32(23);
				b2comp(24) <= B32(24);
				b2comp(25) <= B32(25);
				b2comp(26) <= B32(26);
				b2comp(27) <= B32(27);
				b2comp(28) <= B32(28);
				b2comp(29) <= B32(29);
				b2comp(30) <= B32(30);
				b2comp(31) <= not B32(31);
			elsif (B32(31)='1') then
				b2comp(0) <= B32(0);
				b2comp(1) <= B32(1);
				b2comp(2) <= B32(2);
				b2comp(3) <= B32(3);
				b2comp(4) <= B32(4);
				b2comp(5) <= B32(5);
				b2comp(6) <= B32(6);
				b2comp(7) <= B32(7);
				b2comp(8) <= B32(8);
				b2comp(9) <= B32(9);
				b2comp(10) <= B32(10);
				b2comp(11) <= B32(11);
				b2comp(12) <= B32(12);
				b2comp(13) <= B32(13);
				b2comp(14) <= B32(14);
				b2comp(15) <= B32(15);
				b2comp(16) <= B32(16);
				b2comp(17) <= B32(17);
				b2comp(18) <= B32(18);
				b2comp(19) <= B32(19);
				b2comp(20) <= B32(20);
				b2comp(21) <= B32(21);
				b2comp(22) <= B32(22);
				b2comp(23) <= B32(23);
				b2comp(24) <= B32(24);
				b2comp(25) <= B32(25);
				b2comp(26) <= B32(26);
				b2comp(27) <= B32(27);
				b2comp(28) <= B32(28);
				b2comp(29) <= B32(29);
				b2comp(30) <= B32(30);
				b2comp(31) <= B32(31);
			end if;
			end if;
		end process;
		
		MUX : entity work.two_to_one_mux(behav) port map(B32, b2comp, binvert, bout);
		PASB : entity work.thirty_two_bit_register(behav) port map(bout, clk, rst, pre, ce, output);
end behav;