library IEEE;
use ieee.std_logic_1164.all;

entity d_flip_flop is
	port(
		clk, d, rst, pre, ce : in std_logic;
		q : out std_logic
	);
end d_flip_flop;

architecture behav of d_flip_flop is
begin
	process(clk) is
	begin
		if rising_edge(clk) then
			if (rst='1') then
				q <= '0';
			elsif (pre='1') then
				q <= '1';
			elsif (ce='1') then
				q <= d;
			end if;
		end if;
	end process;
end behav; 
	