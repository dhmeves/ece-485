library IEEE;
use ieee.std_logic_1164.all;

entity multicycle_datapath is
end multicycle_datapath;

architecture behav of multicycle_datapath is

component 