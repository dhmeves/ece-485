library IEEE;
use ieee.std_logic_1164.all;

entity control_unit is
	port(
		op : in std_logic_vector(5 downto 0);
		clk : in std_logic;
		pcWriteCond, pcWrite, IorD, memRead, memWrite, memToReg, irWrite, ALUSrcA, regWrite, regDst : out std_logic;
		pcSource, ALUSrcB, ALUOp : out std_logic_vector(1 downto 0)
	);
end control_unit;

architecture behav of control_unit is
	type states is (S_If, S_Id, S_Ex, S_Mem, S_Wb);
	type operate is (branch, rtype, load, store, jump);
	signal operation : operate;
	signal current_state : states;
	begin
		process(clk) is
		begin
			if rising_edge(clk) then
				if (current_state=S_If) then		
					current_state<=S_Id;
				elsif (current_state=S_Id) then		
					current_state<=S_Ex;
				elsif (current_state=S_Ex) then		
					current_state<=S_Mem;
				elsif (current_state=S_Mem) then		
					current_state<=S_Wb;
				elsif (current_state=S_WB) then	
					current_state<=S_If;
				end if;
			end if;
		end process;
		
		process(current_state) is
		begin
		if (current_state=S_If) then
				pcWriteCond <= '0';
				pcWrite <= '1';
				IorD <= '0';
				memRead <= '1';
				memWrite <= '0';
				memToReg <= '0';
				irWrite <= '1';
				ALUSrcA <= '0';
				regWrite <= '1';
				regDst <= '1';
				pcSource <= "00";
				ALUSrcB <= "01";
				ALUOp <= "00";
			
		end if;

		if (current_state=S_ID) then
				pcWriteCond <= '0';
				pcWrite <= '0';
				IorD <= '0';
				memRead <= '0';
				memWrite <= '0';
				memToReg <= '0';
				irWrite <= '0';
				ALUSrcA <= '0';
				regWrite <= '0';
				regDst <= '0';
				pcSource <= "00";
				ALUSrcB <= "11";
				ALUOp <= "00";
			if (op="000000") then			-- rtype
				operate<=rtype;
			elsif (op="100011") then		-- load
				operate<=load;
			elsif (op="101011") then		-- store
				operate<=store;
			elsif (op="000100") then		-- branch
				operate<=branch;
			elsif (op="010000") then		-- or
				operate<=orop;
			elsif (op="010001") then		-- itype
				operate<=itype;
			end if;
		end if;

		if (current_state=S_Ex) then
				pcWriteCond <= '0';
				pcWrite <= '0';
				IorD <= '0';
				memRead <= '0';
				memWrite <= '0';
				memToReg <= '0';
				irWrite <= '0';
				ALUSrcA <= '0';
				regWrite <= '0';
				regDst <= '0';
				pcSource <= "00";
				ALUSrcB <= "11";
				ALUOp <= "00";
			if (operate=rtype) then			-- add
				--regWrite <= '1';
				--regDst <= '1';
				ALUSrcA <= '1';
				ALUSrcB <= "00";
				ALUOp <= "10";
			elsif (operate=load) then		-- lw
				ALUSrcA <= '1';
				ALUSrcB <= "10";
				ALUOp <= "00";
			elsif (operate=store) then		--sw
				ALUSrcA <= '1';
				ALUSrcB <= "10";
				ALUOp <= "00";
			elsif (operate=branch) then		-- bne/beq
				memToReg <= 'X';
				regDst <= 'X';
				ALUSrcB <= "00";
				ALUOp <= "01";
			elsif (operate=orop) then		-- or
				ALUSrcB <= "00";
				ALUOp <= "00";
			elsif (operate=itype) then		-- andi
				ALUSrcB <= "00";
				ALUOp <= "00";
			end if;
		end if;

		if (current_state=S_Mem) then
			if (op="000000") then			-- add
				pcWriteCond <= '0';
				pcWrite <= '0';
				IorD <= '0';
				memRead <= '0';
				memWrite <= '0';
				memToReg <= '0';
				irWrite <= '0';
				ALUSrcA <= '0';
				regWrite <= '1';
				regDst <= '1';
				pcSource <= "00";
				ALUSrcB <= "00";
				ALUOp <= "10";
			elsif (op="100011") then		-- lw
				pcWriteCond <= '0';
				pcWrite <= '0';
				IorD <= '0';
				memRead <= '1';
				memWrite <= '0';
				memToReg <= '1';
				irWrite <= '0';
				ALUSrcA <= '1';
				regWrite <= '1';
				regDst <= '0';
				pcSource <= "00";
				ALUSrcB <= "00";
				ALUOp <= "00";
			elsif (op="101011") then		--sw
				pcWriteCond <= '0';
				pcWrite <= '0';
				IorD <= '0';
				memRead <= '0';
				memWrite <= '1';
				memToReg <= 'X';
				irWrite <= '0';
				ALUSrcA <= '1';
				regWrite <= '0';
				regDst <= 'X';
				pcSource <= "00";
				ALUSrcB <= "00";
				ALUOp <= "00";
			elsif (op="000100") then		-- bne/beq
				pcWriteCond <= '0';
				pcWrite <= '0';
				IorD <= '0';
				memRead <= '0';
				memWrite <= '0';
				memToReg <= 'X';
				irWrite <= '0';
				ALUSrcA <= '0';
				regWrite <= '0';
				regDst <= 'X';
				pcSource <= "00";
				ALUSrcB <= "00";
				ALUOp <= "01";
			elsif (op="010000") then		-- or
				pcWriteCond <= '0';
				pcWrite <= '0';
				IorD <= '0';
				memRead <= '0';
				memWrite <= '0';
				memToReg <= '0';
				irWrite <= '0';
				ALUSrcA <= '0';
				regWrite <= '0';
				regDst <= '0';
				pcSource <= "00";
				ALUSrcB <= "00";
				ALUOp <= "00";
			elsif (op="010001") then		-- andi
				pcWriteCond <= '0';
				pcWrite <= '0';
				IorD <= '0';
				memRead <= '0';
				memWrite <= '0';
				memToReg <= '0';
				irWrite <= '0';
				ALUSrcA <= '0';
				regWrite <= '0';
				regDst <= '0';
				pcSource <= "00";
				ALUSrcB <= "00";
				ALUOp <= "00";
			end if;	
		end if;

		if (current_state=S_Wb) then
			if (op="000000") then			-- add
				pcWriteCond <= '0';
				pcWrite <= '0';
				IorD <= '0';
				memRead <= '0';
				memWrite <= '0';
				memToReg <= '0';
				irWrite <= '0';
				ALUSrcA <= '0';
				regWrite <= '1';
				regDst <= '1';
				pcSource <= "00";
				ALUSrcB <= "00";
				ALUOp <= "10";
			elsif (op="100011") then		-- lw
				pcWriteCond <= '0';
				pcWrite <= '0';
				IorD <= '0';
				memRead <= '1';
				memWrite <= '0';
				memToReg <= '1';
				irWrite <= '0';
				ALUSrcA <= '1';
				regWrite <= '1';
				regDst <= '0';
				pcSource <= "00";
				ALUSrcB <= "00";
				ALUOp <= "00";
			elsif (op="101011") then		--sw
				pcWriteCond <= '0';
				pcWrite <= '0';
				IorD <= '0';
				memRead <= '0';
				memWrite <= '1';
				memToReg <= 'X';
				irWrite <= '0';
				ALUSrcA <= '1';
				regWrite <= '0';
				regDst <= 'X';
				pcSource <= "00";
				ALUSrcB <= "00";
				ALUOp <= "00";
			elsif (op="000100") then		-- bne/beq
				pcWriteCond <= '0';
				pcWrite <= '0';
				IorD <= '0';
				memRead <= '0';
				memWrite <= '0';
				memToReg <= 'X';
				irWrite <= '0';
				ALUSrcA <= '0';
				regWrite <= '0';
				regDst <= 'X';
				pcSource <= "00";
				ALUSrcB <= "00";
				ALUOp <= "01";
			elsif (op="010000") then		-- or
				pcWriteCond <= '0';
				pcWrite <= '0';
				IorD <= '0';
				memRead <= '0';
				memWrite <= '0';
				memToReg <= '0';
				irWrite <= '0';
				ALUSrcA <= '0';
				regWrite <= '0';
				regDst <= '0';
				pcSource <= "00";
				ALUSrcB <= "00";
				ALUOp <= "00";
			elsif (op="010001") then		-- andi
				pcWriteCond <= '0';
				pcWrite <= '0';
				IorD <= '0';
				memRead <= '0';
				memWrite <= '0';
				memToReg <= '0';
				irWrite <= '0';
				ALUSrcA <= '0';
				regWrite <= '0';
				regDst <= '0';
				pcSource <= "00";
				ALUSrcB <= "00";
				ALUOp <= "00";
			end if;
		end if;
	end process;
end behav;